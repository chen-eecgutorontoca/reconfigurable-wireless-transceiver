

module tx_vga(
    input logic clk,
    input logic rst_n,
    output logic tx_vga_sclk,
    output logic tx_vga_CS,
    output logic tx_vga_SDO,
    input logic tx_vga_SDI
);



